BZh91AY&SY=�j� �߀Py���߰����`�8�ˤ��ڪxE
 A(�5<�L!4��2m@ �  ��M�(��h ��@�j&��( dd=@    S����� �d�L��M4  ���a2dɑ��4�# C T��=L���6��HGꌁ����3SH8v���3I!�~4Ē��՟��eH��H��Q�~�Uǻ)#Ip�Z�"K�z�Ic�/���xߩ��          @ A�  @       ��   %���Q�Z���UM_��W,��=:��]��囪���q��GnEC�6ݫmY�e�}�Z�R�[*�n�Uʱ�4�SiVf6Uj�>x&�1!26��nZ`@Z(�N8�s�u�!u� @)��Ҟ<���:[R۞�=`  b�  4� (@  �  ؀    c�]����	&�M?>��t!�n�1��C��gae��LΈ�1:�� �֦�)��*�����E�){^T�\�8S��R�)��n�8O�*���a$�o�k�OIt�P 1&�wK�.���7�D�!�+��Z���։WR�Fw�`o���"),��S�˺����T�$kWZ;kI(��]��L���~��0  ���$�T�*u��niuǇN�1�I�m�Jک�Ҕ��K�K��2�q�*th�6�]��8�7ɘ}q������[��  4��}��[T�f��m.SN�K8�Q.]�/��k+[�x��"�啔T��Y=�B'�i%�bk:�֪7Ǣ��|�  ^m�[l���@�JBq����Lۙ�[��EΚ���E6���ee��m������Ko*.��Vs�n�.�y���x�zAtk��Z��y��K�a�\�ɩ��k{�rqj���v��h
2�:B}P <2���/C�D�V��E����sf���A\�\"�I��el�V��X  WI����^�7��g��Ҭ��!m��4�޵���k3s���r��Gx��wO׵�  h����͕��b�ۨ�����TF#��u�k:�&mGCqɵ�d.  Z�w���3C=J��,U5����Pdq�+{�Y�F^��y�7wd�2K�U*�$����|���f�&L�Ҽ�{3b�C5(�)eK�*QE(�ER�LQR��R��S�e�*���b�j*QJ)E*Q��֒gQ�E��U�KYe��{�`�u����L����n"J�!U-������S��4��S2��I+4��Ij/�.��mQ�{ )�۽�rF%y�ѣ+�aX"�+���<u���M��"
�
�Ϣow�9�#w�^�q���OG�Tē���#T�;���{=�FjQ}:[*��ձ%c&:�tK�6���PT�nj�U%m�X**��"�@�P[.ԥ�Η������I�z[�ە��R�AV�������e��̮��J�U��`͇����xgǌ��_%�L������}��u�h��Q��^5� R\X8h�kA�I%+h�@7�*��?8͊�э9���\$9ȃ�}{L��͏
z�,��[���a�LIߖ]IL�aǥ���u,���~yKgӻ&v���si�*x���.�4y3��E/��y;dW_���;,�wK|�>>�����X��7..�|�,}xF�;�f�
�'qJ>__�DOOnn��7m,�w`�|gTm-����1��V�>ku�������MX5��t��F�1�vR κxn��y���t)���K��/f��>V�jШ��4:��b	?N2f�'���S���� �u��P1((�ȗ��.�p� {��|