BZh91AY&SYH�� �_�Py���߰����`�8z��Ӥ����B@@I"d�ѩ&�ީ���4y@�4 i���	�$��#@ �  ��&RP�`�	� 	��	4       9�14L�2da0M4����DF�{(�2�Sѩ���   3$���Db$D�$���hC2K��?�#J����VT���.#Ӥ��YM-����=��,=���^r�z:}*�  0�         @  �   @      �.W����k�ǲ�|��f�G�B
|���F8f�lF�fk5��R�����Pꋷef�%�Z(K��{����������JU�J��Hf��s�͟��^�+O�T��F���d���lE�"2x�^��yO?/��]7���I�Ͷ�i��{a�[m��n�p�n[m�e��m��m�e��vۆ�a��m��l6�m�e�]xy��� ��R=B��T
��IGx�"8t�`�$L# F��ZI$��Cv(+���Mn�dQ��X,stP��[6?[9�p�瞁�@�ûZ �U�Ϳ��K}�  @�I�_Ĵ�q;S�ҍ��25��Z�jm@�p2�q���L�"�a�Z֤�q�ʗšӨ�G8��--�IEO�������7�`  �k�	��*u��Zl�a��{�:�wa.@ì����
��:eVVr��� 8pb�D����xk]�"   6Vz|3�T�b��WKI�A��e� ��Wh�'r.�v
�HaU��XACf�!B@� l�7�L�TR%�b�   
�.ݕ�%�� p�	���A{1F�֞+"�*RI7�I��j�3�}�|�Wx��"�KZ-@ s	MM='.���{3J�3d�Nȓi�K�cXѭLV3���S��P�A*	�OI$ID�wS-D��&z�c�=]�s�sjy�W|�#-*������f�I$��E]7e,�UL�w'dQ��ȼ#a��A53NPo��Q�������Q2�3��RI$�FE<����ӥ�V0�%��=����n_"D;|�Qv��JI$���U8��HWhnv(Ps��(���iB�-�e����r7�^��� �A����a����{�I���VZ3��3�5�����e.��f.)JYK)JV.̌JYK)T�����KKK.j0���U*�F0Fړ[41���,�R��Y��^[��1Z���v"KdC2��w:��z]�Q�%^6�����>���C�d9G3��Pp>�������=a)������xP�8�u;���1�e�I��dA�Ƀޜ�۞:hn�eVb?����}r��>	���6��ۇ�������U�:6��6�\��Lj�Dw�g��0�oҧ��b/�\��j�I�6H7*��J�3kc���7I�y�����e�����M����|�j^�_����i2j˽�I��k�|�dA�ج�w�����}^~7����)�(��z[��eG��Q�(d�� <VfE٩Hj�%4E�&�	���nI��.�<������76̵��2v駉+No�h$)��j��1�I���eq����5��vY�V.�1��bA�Ьu��\����"�{A��昧�ݮ���Ns���w�R����FX�^�,ۡ �d�*�ߣ�"盯W?�ɳw)�h�ɯ4ki�a��d���C����kg�O��NFM��N�_���[RB�����`6��լd:���V�!h�u�Gk�_Ǥqe���hV�F#����릗3ATz�r��"Eƹ�ܑN$.4�@