BZh91AY&SY�� ,_�Px��g߰����  `�<o�(���B��_�MM�#Sz��j�h�2hP 50hҔԀM  d�  T�CA%M��@�  h  	O�H����4`	�&C��F&�	�&�`�i���!��!��$�jz���i� i�Q5 3�BH 4B�@$�o���8���{���$�d��u��vM$��,��2�5f��q-�r3�s�n_�W(  @     � ��mm��~����x�M����{I�\OR����-��P��e�+.��;�TS�ɶ���N��E� ͛��m�NQqA��-
ʊW�ڦ'?K��N� �� H~X�˂��p��[��)�,�4� ��R@.|���zf�=���%	$�I:I$��I$�I$�Wwwe�X�$�Ibd�I�$���T�P�K3.��=��w����9������Be�逿AW	��l�P�*�Kﺔ�)J�o����a%��('����.�l��bna�����  0��5ldP<� ��8I$�$'x�����XCrUT�Q���y�ߕ�r1�!� �����ĵ�Q6�嵰�<��~��9��8䨙��I$�����P[u!KJ`�;�ⴟJ*.�܆f�5�.���ᦃ�wDL�i
�gQ����otn:���W��I'�!�Cddū7dPM-m��<�s{S�:�����񓖶��E�l���P������M���`9Y8�$�q,���i0_�.��8*���ne����&yy�+!�E�Cҁ��D7X]ZT�о�cgj������h����y��J���d�� ��z�(��@aa�1�!�M�i$��U)��!�ҙ;:���X�����!�D�C[�� �MS�$�����I%��6���]<n���&-H�ڗa��Bx�3���C�f���:;c�ު���&y��#���J�k=9]��ˮ�Ya��D��?[OH�j{buo�MIx�I!^憡Z7PV�Z�)��2������������H �O����w<��j�n�\-���r��>�͕������Rg�j�$���Ĥ�Jl�X�������bV�V�����$�5�ij����֪2Ii��Z��[�4�6��C*km�� I�&�W�u#��<�)������j�z�|~��ċ�h�z{n���b{���I�>P�-,  ��0���?r�z�X������'��Ѩ,���I�����ܪ�����0�������jU&5k2.{�G�%��ȥ+��C���ie����C\\�JƁ����PO�Lj�!����KJ�;A!��!��F��uZ�K�YA����L���\�{v�e�*��$�M�sc�����u&�3�ͤ��H��L�2��g�Zb�In�Ų1V���Xr0�D
�J����nN-���\���D�B�W���2W)�"b-d8�@L�I8��(dR���_9r��7�  ��29zz5�zs�I+��㤱��n@��՝���#ã����H���q���� �#jc[7�I$��)*�!kF�*X�6�A��@�(��Ȩ�%�]zZمvzi�!:L�YR��2��)�9�.�f(쮰�S�&d�ܢ��Ae�i�ĮnS	%��'~��{J�3!q��3h�>`��H�
� 1�