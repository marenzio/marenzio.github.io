BZh91AY&SY�1�j $߀Pxg��g߰����`n��� ���Z��(�=4'�l����aSA��MPz@�ƃJP��hC@  ��T����Ѡ�M�A�LC@ 	4����P�hh=L�   hP4d���`F�b0L�`�M	��zdi4�)���F� h z�E�b�J�%@�Xk�Q���������&��Y��ރ�Ȅ&����r�O
f�q�=�f�͊�������������������������6op7#�a���n%d�`��0c ��b�V����aL�z���Ȇ1F�Q�艆ɖ�Rb�$�d�f�N	���>n|3k�I��#d�Q�^V��u
�'�D�	֙D@^�-����������K����������$�I$�JRH��I,�̬�С�I%i$�V���I$�t�K����;�pq�q�7���<C�g=���U�j�
���a$�P�<�DK�f��"X��W�,|�R�Y�r-���%E^Eev�ps�s(�#�`&{%L���H��f �/�Dv�����ʇ�nS	};0���Y����	?)��~�氆�r�v����2�ٽ9f��ro��&fdI�:�<�yu�� cph�ql3\>>�%�)�ȶ�&Z1���(~u�PE�x�0�Q�Lɞ8b�Q�h��a�:��qp��o���L���0��S�`���r�A��1
a�d�I�`S;U�T@�����5Ĉ��N@��!���H�D��Ql40Y=�)]N
R�I$�
����v	�H{����r��f�y���wl�l�,�I��I˚�E�C�]cu�ȘWq�P֍"�2x`���� [ޒI+\�Nضt��(�<�l6�7Y�n�/mǔ��:��M�uղȗ7y���3�W]�p��Bf�����h����EբI.A��&^�v�,�WR猘�V�z{��ꎼ�<����%T����l���]F0a��^�B"&�YZ""1�FW<���Ds�����$�F#U
"1��"`�b"1���%-�+��mLFW��r�ML��w��D
���T���dW�Ã.>��M;��U�o�}FrJ��ɼ�|����8�8�}he.'z�-���tu���S9�7����w��k��6Ӵp�#�� d<���Y��]�p�lшe6�_� ��(#֕�Q�S@x?�C̡�׎�}�&x��8֑+L��(����A��8�2��!\�$�i��&[�Fk���X��<�&�Y�4�����L�C�$_.���,��#I1��"�0�=#��U��A��L�㛓��6��Qm��!�Ƞv��QR�dJf݄�_�+�%�\Z�:q6�y`F�\De���ka��]��3�w���S���D��xZL�I���w�{����A	0Z�]m� }d�N��_u�@n��,ӀJ�C;Y��5HBP�1�]{D6�Y�B�[��� ���}�����&s5��<����rЎC�ɉ��">3zF��-��!bܶ8�;m7:� �TD� ���c�T��p֤�I��o���5N<%|ǐE=��)56'��n)p\2u62,J�@子	�GA}ᗤ�m�0�n,zAm:�z5\̲Q�Ɔ�Kk ����.�p�!�cB�