BZh91AY&SY�<hA �_�Pxg��g߰����`�����` �^I�&����MOM!��� h24���i*% �`�	�` �j���zI� 0   &j�H�S�1�=5  20��@mT�h@�4    ��S�i52bi���  �dd��@��	4!��C(�h'���
�-� �l'� ���ZV�{�y֤�%��t�� � �  �  [w«�������-LQ�ӋN��}}��6�ʙ�,��L�>+.�D,^���qՋ7B�4�
��l��oUp�R��G5�b1�F��#���f�AB������Z�2[e��-��rt�I$�I$���$�$��$���$�I%)$�I)I:Jd��?�_8 ��.����5������=�J,�rsV���\�$��S33F9(p}��F��~ ǚo�1���Iyhg��C��+0���9�8���}��0�J��I%��p&
�g���Ty;�bX��f�h�T&�#&�
-�ІN�x���f?e�"I'���ޚ�=��jh`̱ݰ��9��Xm/�kg��,7��VPвoZ7��3�=$��l]�l�79��a�����O��O�mLT4J�bnC��I6�<�zV�+�2�p4�ˇ�n��fʥ����r�0N5�(Oc�Z�0�TEÂ,�xgb���#5����{~�d�=kg�"���WT8Fc���HR1a�н�\����s��:���I(�G�T\��*��u�̫x.&i�*�·���;��H��-ڥ���^QΩ�ϡ��`���ˎ�SiM��/3�	��S��ܕ;��d]�"T4Z�����3�* ;)�q0#��\�U�^�A��-%�T��������+{˸j����F�sM�7V%��RY �D� ��	!$$�U$$������lL���<�s^�5���́�T���[���1�̌���wJk���~o�-B��2�?;����h�����vY�[?�?��M�����.������<��(�� ��	��T���k���J^��9%���0�,� ���f
#�LY��\4�h����G�5��Нu�8P��ӋB��ᤲ7�OC]�D+1	Y�`&S|Lj�s!�Z�|�9��m�v�����u&u�s�U�f��Ø�#D�<%��ߺؘ ��9��m���SF��@�d�h�4����g���@�b�B"Z�Ā[�,f�o;�V�~��Q��B� iu���Gkr�X*Ma9)��
����SD�Ba� .�}�H�r����}Q �b��g �sX��t�!��28��8=�[� ��s�R�ܴ�z��8Tt8�����nP��@�6�i�u,��6��I�X�0H�6i���2�8�21z�Q�!`kȐ��4P<MZ�u\�n��Z���ו��M�BpƉ �w����b��J�7����ˈ��@砪���q=(+��L���5׽v_K2�I/�&�KAp��]��BC��